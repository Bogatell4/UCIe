
module LTSM_top (

    input clk_100MHz,
    input reset,
    input enable_i,

    input MB_

    
);




end module;
